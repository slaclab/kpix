-------------------------------------------------------------------------------
-- Title      : Standard RTL Package
-------------------------------------------------------------------------------
-- File       : StdRtlPkg.vhd
-- Author     : Benjamin Reese 
-- Standard   : VHDL'93/02, Math Packages
-------------------------------------------------------------------------------
-- Description: This package defines "sl" and "slv" shorthand subtypes for
--              std_logic and std_logic_vector repectively.  It also defines
--              many handy untility functions. Nearly every .vhd file should
--              use this package.
-------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

package StdRtlPkg is

  -- Typing std_logic(_vector) is annoying
  subtype sl is std_logic;
  subtype slv is std_logic_vector;

  -- Very useful functions
  function log2(constant number : integer) return integer;
  function bitReverse (a         : slv) return slv;

  -- This should be unnecessary in VHDL 2008
  function toBoolean (logic : sl) return boolean;
  function toSl (bool       : boolean) return sl;

  -- Unary reduction operators
  function uOr (vec      : slv) return sl;
  function uAnd (vec     : slv) return sl;
  function uXor (vec     : slv) return sl;
  function uOrBool (vec  : slv) return boolean;
  function uAndBool (vec : slv) return boolean;
  function uXorBool (vec : slv) return boolean;

  -- Avoid bla = "00000" literal comarisons that don't scale naturally with bla'length
  function slvZero (length      : integer) return slv;
  function unsignedZero (length : integer) return unsigned;
  function isZero (vec          : slv) return boolean;
  function isZero (vec          : unsigned) return boolean;

  -- Create an slv of given size with every v
  function slvAll (value : sl; length : natural) return slv;

  -- These just use uXor to calulate parity
  -- Output is parity bit value needed to achieve that parity given vec.
  function evenParity (vec : slv) return sl;
  function oddParity (vec  : slv) return sl;

  -- Gray Code functions
  function grayEncode (vec : unsigned) return unsigned;
  function grayEncode (vec : slv) return slv;
  function grayDecode (vec : unsigned) return unsigned;
  function grayDecode (vec : slv) return slv;


  -- Some synthesis tools wont accept unit types
  --type frequency is range 0 to 2147483647
  --  units
  --    Hz;
  --    kHz = 1000 Hz;
  --    MHz = 1000 kHz;
  --    GHz = 1000 MHz;
  --  end units;

  --function toTime(f : frequency) return time;

end StdRtlPkg;

package body StdRtlPkg is


  ---------------------------------------------------------------------------------------------------------------------
  -- Function: log2
  -- Purpose: Finds the log base 2 of an integer
  -- Input is rounded up to nearest power of two.
  -- Therefore log2(5) = log2(8) = 3.
  -- Arg: number - integer to find log2 of
  -- Returns: Integer containing log base two of input.
  ---------------------------------------------------------------------------------------------------------------------
  function log2(
    constant number : integer)
    return integer
  is
    variable divVar : integer;
    variable retVar : integer := 0;
  begin
    divVar := number;

    while (divVar /= 1) loop
      if (divVar mod 2 > 0) then
        retVar := retVar + 1;
      end if;
      divVar := divVar/2;
      retVar := retVar + 1;
    end loop;
    return retVar;
  end function log2;

  function bitReverse (a : slv)
    return slv
  is
    variable resultVar : slv(a'range);
    alias aa           : slv(a'reverse_range) is a;
  begin
    for i in aa'range loop
      resultVar(i) := aa(i);
    end loop;
    return resultVar;
  end;

  function toBoolean (
    logic : sl)
    return boolean is
  begin  -- function toBoolean
    return logic = '1';
  end function toBoolean;

  function toSl (
    bool : boolean)
    return sl is
  begin  -- function toSl
    if (bool) then
      return '1';
    else
      return '0';
    end if;
  end function toSl;

  ---------------------------------------------------------------------------------------------------------------------
  -- Unary reduction operators
  ---------------------------------------------------------------------------------------------------------------------
  function uOr (vec : slv) return sl is
  begin
    for i in vec'range loop
      if (vec(i) = '1') then
        return '1';
      end if;
    end loop;
    return '0';
  end function uOr;

  function uAnd (vec : slv) return sl is
  begin
    for i in vec'range loop
      if (vec(i) = '0') then
        return '0';
      end if;
    end loop;
    return '1';
  end function uAnd;

  function uXor (vec : slv) return sl is
    variable intVar : sl;
  begin
    for i in vec'range loop
      if (i = vec'left) then
        intVar := vec(i);
      else
        intVar := intVar xor vec(i);
      end if;
    end loop;
    return intVar;
  end function uXor;

  function uOrBool (vec : slv) return boolean is
  begin
    return toBoolean(uOr(vec));
  end function;

  function uAndBool (vec : slv) return boolean is
  begin
    return toBoolean(uAnd(vec));
  end function;

  function uXorBool (vec : slv) return boolean is
    variable intVar : sl;
  begin
    return toBoolean(uXor(vec));
  end function;

  ---------------------------------------------------------------------------------------------------------------------
  -- Functions to get a vector of all same value
  ---------------------------------------------------------------------------------------------------------------------
  function slvAll (value : sl; length : natural) return slv is
    variable retVar : slv(length-1 downto 0) := (others => value);
  begin
    return retVar;
  end function;

  function slvZero (length : integer) return slv is
  begin
    return slvAll('0', length);
  end function;

  function unsignedZero (length : integer) return unsigned is
  begin
    return unsigned(slvZero(length));
  end function;

  function isAll (vec : slv; value : sl)
    return boolean is
  begin
    return vec = slvAll(value, vec'length);
  end function;

  function isZero (vec : slv)
    return boolean is
  begin
    return vec = slvZero(vec'length);
  end function;

  function isZero (vec : unsigned)
    return boolean is
  begin
    return vec = unsignedZero(vec'length);
  end function;




  -----------------------------------------------------------------------------
  -- Functions to determine parity of arbitrary sized slv
  -----------------------------------------------------------------------------
  -- returns '1' if vec has even parity
  function evenParity (vec : slv)
    return sl is
  begin
    return not uXor(vec);
  end function;

  -- return '1' if vec has odd parity
  function oddParity (vec : slv)
    return sl is
  begin
    return uXor(vec);
  end function;

  -----------------------------------------------------------------------------
  -- Functions for encoding and decoding grey codes
  -----------------------------------------------------------------------------
  -- Get next gray code given binary vector
  function grayEncode (vec : unsigned)
    return unsigned is
  begin
    return vec xor shift_right(vec, 1);
  end function;

  -- SLV variant
  function grayEncode (vec : slv)
    return slv is
  begin
    return slv(grayEncode(unsigned(vec)));
  end function;

  -- Get the binary equivalent of a gray code created with gray_encode.
  function grayDecode (vec : unsigned)
    return unsigned is
    variable retVar : unsigned(vec'range) := (others => '0');
  begin
    for i in vec'range loop
      if (i = vec'left) then
        retVar(i) := vec(i);
      else
        if (vec'ascending) then
          retVar(i) := retVar(i-1) xor vec(i);
        else
          retVar(i) := retVar(i+1) xor vec(i);
        end if;
      end if;
    end loop;
    return retVar;
  end function;

  -- SLV variant
  function grayDecode (vec : slv)
    return slv is
    variable retVar : slv(vec'range) := (others => '0');
  begin
    return slv(grayDecode(unsigned(vec)));
  end function;

  ---------------------------------------------------------------------------------------------------------------------
  -- Convert a frequency to a period (time).
  ---------------------------------------------------------------------------------------------------------------------
  --function toTime(f : frequency) return time is
  --begin
  --  return(1.0 sec / (f/Hz));
  --end function;
  
end package body StdRtlPkg;
